module fpu_64_divider_tb ();
    
    parameter WIDTH = 64;
    reg [WIDTH-1:0] A;
    reg [WIDTH-1:0] B;
    wire [WIDTH-1:0] result;
    wire overflow;
    wire underflow;

    fpu_64_divider #(.WIDTH(WIDTH)) uut (
        .A(A),
        .B(B),
        .result(result),
        .overflow(overflow),
        .underflow(underflow)
    );

    initial begin
        $monitor("A = %h | B = %h | Result = %h | Overflow = %b | Underflow = %b", A, B, result, overflow, underflow);
        // Test case 1: 4.0 / 2.0
        A = 64'b0100000000010000000000000000000000000000000000000000000000000000; // 4.0
        B = 64'b0100000000000000000000000000000000000000000000000000000000000000; // 2.0
        #10;

        // Test case 2: 1.0 / 0.5
        A = 64'b0011111111110000000000000000000000000000000000000000000000000000; // 1.0
        B = 64'b0011111111100000000000000000000000000000000000000000000000000000; // 0.5
        #10;

        // Test case 3: 2.0 / 4.0
        A = 64'b0100000000000000000000000000000000000000000000000000000000000000; // 2.0
        B = 64'b0100000000010000000000000000000000000000000000000000000000000000; // 4.0
        #10;

        // Test case 4: Division by zero (B=0)
        A = 64'b0100000000000000000000000000000000000000000000000000000000000000; // 2.0
        B = 64'b0000000000000000000000000000000000000000000000000000000000000000; // 0.0
        #10;

        // Test case 5: Zero divided by a number (A=0)
        A = 64'b0000000000000000000000000000000000000000000000000000000000000000; // 0.0
        B = 64'b0100000000000000000000000000000000000000000000000000000000000000; // 2.0
        #10;
        
        $finish();
    end
endmodule